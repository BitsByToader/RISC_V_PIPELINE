`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/11/2023 08:58:41 PM
// Design Name: 
// Module Name: instruction_decode
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instruction_decode(
    input clk,
    input reset,
    input flush_pipe,

    // From Hazard Detection Unit
    input stall_pipeline,

    // from IF
    input [31:0] pc_addr_in,
    input [31:0] instr,
    
    // From WB
    input [4:0] write_reg_wb,
    input [31:0] data_reg_wb,
    input regwrite_ctrl_wb,
    
    // Pipeline reg ID->EX
    output reg [31:0] pc_addr_out,
    output reg [31:0] rd1,
    output reg [31:0] rd2,
    output reg [31:0] imm_gen_out,
    output reg [6:0] funct7,
    output reg [2:0] funct3,
    output reg [4:0] write_reg_out, // or rd
    output reg [4:0] rs1_out,
    output reg [4:0] rs2_out,
    
    // Output from Control Module
    output reg mem_read_ctrl,
    output reg mem_write_ctrl,
    output reg mem_to_reg_ctrl,
    output reg reg_write_ctrl,
    output reg branch_ctrl,
    output reg unconditional_branch_ctrl,
    output reg alusrc_a_ctrl,
    output reg [1:0] alusrc_b_ctrl,
    output reg addr_src_ctrl,
    output reg [1:0] aluop_ctrl
);

    // Generated by the regfile
    wire [31:0] rd1_tmp; // ~~ reg data 1 
    wire [31:0] rd2_tmp; // ~~ reg data 2
    
    // Generated by the imm gen
    wire [31:0] imm_gen_out_tmp;
    
    // Generated by the control module
    wire mem_read_ctrl_tmp;
    wire mem_write_ctrl_tmp;
    wire mem_to_reg_ctrl_tmp;
    wire reg_write_ctrl_tmp;
    wire branch_ctrl_tmp;
    wire unconditional_branch_ctrl_tmp; // For jump instructions!
    wire alusrc_a_ctrl_tmp; // For jump instruction!
    wire [1:0] alusrc_b_ctrl_tmp; // For jump instruction!
    wire addr_src_ctrl_tmp; // For jumps!
    wire [1:0] aluop_ctrl_tmp;

    register_file regfile(
        .clk(clk),
        .reset(reset),
        .wen(regwrite_ctrl_wb),
        .ra(instr[19:15]),
        .rb(instr[24:20]),
        .rc(write_reg_wb),
        .da(rd1_tmp),
        .db(rd2_tmp),
        .dc(data_reg_wb)
    );
    
    imm_gen immgen(
        .instr(instr),
        .imm(imm_gen_out_tmp)
    );
    
    // From here on out I got too bored to write the module instantiation like above :-)
    // Even though it might lead to my demise :-)
    control_module ctrl(
        instr[6:0],
        stall_pipeline,
        mem_read_ctrl_tmp,
        mem_to_reg_ctrl_tmp,
        mem_write_ctrl_tmp,
        reg_write_ctrl_tmp,
        branch_ctrl_tmp,
        unconditional_branch_ctrl_tmp, // For jump instructions!!
        alusrc_a_ctrl_tmp, // For jump instructions!
        alusrc_b_ctrl_tmp,  // For jump instructions!
        addr_src_ctrl_tmp, // For jumps!
        aluop_ctrl_tmp
    );
    
    // Pipeline registers
    always @(posedge clk) begin
        if ( reset || flush_pipe ) begin
            pc_addr_out <= 0;
            rd1 <= 0;
            rd2 <= 0;
            imm_gen_out <= 0;
            funct7 <= 0;
            funct3 <= 0;
            write_reg_out <= 0;
            rs1_out <= 0;
            rs2_out <= 0;
            mem_read_ctrl <= 0;
            mem_write_ctrl <= 0;
            mem_to_reg_ctrl <= 0;
            reg_write_ctrl <= 0;
            branch_ctrl <= 0;
            unconditional_branch_ctrl <= 0; // For jumps!
            alusrc_a_ctrl <= 0; // For jumps!
            alusrc_b_ctrl <= 0; // For jumps!
            addr_src_ctrl <= 0;
            aluop_ctrl <= 0;
        end else begin
            pc_addr_out <= pc_addr_in;
            rd1 <= rd1_tmp;
            rd2 <= rd2_tmp;
            imm_gen_out <= imm_gen_out_tmp;
            funct7 <= instr[31:25];
            funct3 <= instr[14:12];
            write_reg_out <= instr[11:7];
            rs1_out <= instr[19:15];
            rs2_out <= instr[24:20];
            mem_read_ctrl <= mem_read_ctrl_tmp;
            mem_write_ctrl <= mem_write_ctrl_tmp;
            mem_to_reg_ctrl <= mem_to_reg_ctrl_tmp;
            reg_write_ctrl <= reg_write_ctrl_tmp;
            branch_ctrl <= branch_ctrl_tmp;
            unconditional_branch_ctrl <= unconditional_branch_ctrl_tmp; // For jumps!
            alusrc_a_ctrl <= alusrc_a_ctrl_tmp; // For jumps!
            alusrc_b_ctrl <= alusrc_b_ctrl_tmp; // For jumps!
            addr_src_ctrl <= addr_src_ctrl_tmp; // For jumps!
            aluop_ctrl <= aluop_ctrl_tmp;
        end
    end
    
endmodule